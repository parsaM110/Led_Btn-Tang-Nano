module led_btn(
    input btn_i,
    output led_o
);

assign led_o = btn_i;

endmodule